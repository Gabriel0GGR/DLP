-- Contador de decada sincrono "UP/DOWN"
-- Exemplo em VHDL

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity contador_ud is
	port
	(
		clk, reset, ud, enable: in std_logic;
		Q0, Q1, Q2, Q3, CY: out std_logic
	);
end contador_ud;

architecture comportamento of contador_ud is

	signal cont: unsigned(3 downto 0);

begin
	process(clk, reset, ud) is
	begin
		if reset='0' then cont<="0000";
		elsif clk'event and clk='0' and enable='1' then
			if ud='1' then
				if cont="1001" then cont<="0000";
					CY<='0';
				else cont<=cont+1;
					CY<='1';
				end if;
			else
				if cont="0000" then cont<="1001";
					CY<='0';
				else cont<=cont-1;
					CY<='1';
				end if;
			end if;
		end if;
	end process;
	
	Q0<=cont(0);
	Q1<=cont(1);
	Q2<=cont(2);
	Q3<=cont(3);
	
end comportamento;